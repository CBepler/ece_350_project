module or32(Out, A, B);
    
    input [31:0] A, B;
    output [31:0] Out;

    or or0(Out[0], A[0], B[0]);
    or or1(Out[1], A[1], B[1]);
    or or2(Out[2], A[2], B[2]);
    or or3(Out[3], A[3], B[3]);
    or or4(Out[4], A[4], B[4]);
    or or5(Out[5], A[5], B[5]);
    or or6(Out[6], A[6], B[6]);
    or or7(Out[7], A[7], B[7]);
    or or8(Out[8], A[8], B[8]);
    or or9(Out[9], A[9], B[9]);
    or or10(Out[10], A[10], B[10]);
    or or11(Out[11], A[11], B[11]);
    or or12(Out[12], A[12], B[12]);
    or or13(Out[13], A[13], B[13]);
    or or14(Out[14], A[14], B[14]);
    or or15(Out[15], A[15], B[15]);
    or or16(Out[16], A[16], B[16]);
    or or17(Out[17], A[17], B[17]);
    or or18(Out[18], A[18], B[18]);
    or or19(Out[19], A[19], B[19]);
    or or20(Out[20], A[20], B[20]);
    or or21(Out[21], A[21], B[21]);
    or or22(Out[22], A[22], B[22]);
    or or23(Out[23], A[23], B[23]);
    or or24(Out[24], A[24], B[24]);
    or or25(Out[25], A[25], B[25]);
    or or26(Out[26], A[26], B[26]);
    or or27(Out[27], A[27], B[27]);
    or or28(Out[28], A[28], B[28]);
    or or29(Out[29], A[29], B[29]);
    or or30(Out[30], A[30], B[30]);
    or or31(Out[31], A[31], B[31]);
    
endmodule
